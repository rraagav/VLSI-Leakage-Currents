*CONDUCTION NMOS W1

.INCLUDE 45nm_MGK.pm
.OPTIONS GMIN=1e-020 ABSTOL=1e-18 TEMP=85

*Definizione dei parametri
.PARAM Lmin=45n
.PARAM Wmin=90n
.PARAM Ldiff=45n
.PARAM supply=1.1


.GLOBAL gnd

M1 drain1 gate1 net1 body1 nmos W={Wmin} L={Lmin} AS={Wmin*Ldiff} AD={Wmin*Ldiff} PS={2*(Ldiff+Wmin)} PD={2*(Ldiff+Wmin)}
M2 net2  gate2 source2 body2 nmos W={Wmin} L={Lmin} AS={Wmin*Ldiff} AD={Wmin*Ldiff} PS={2*(Ldiff+Wmin)} PD={2*(Ldiff+Wmin)}

*NMOS Turned on
Vd drain1 gnd 1.1
Vg1 gate1 gnd 0
Vg2 gate2 gnd 0
Vb1 body1 gnd 0
Vb2 body2 gnd 0
Vs2 source2 gnd 0
Vd2 net1 net2 0
*Vdd alim 0 0


.CONTROL
*let voltage=0
*let Vddbasic=1.1
*while voltage le Vddbasic
*  let voltage = voltage + 0.05
*  alter sw = voltage
dc Vd 0 1.1 0.05
echo V(drain1) V(gate1) V(net1) V(body1) I(Vd) I(Vg1) I(Vd2) I(Vb1) V(net2) V(gate2) V(net2) V(body2) I(Vd2) I(Vg2) I(Vs2) I(Vb2)  > NMOS_Stack_00_W1.txt
let i=1
while (i <= length(V(drain1)))
    let Vdrain1 = V(drain1)[i]
    let Vgate1 = V(gate1)[i]
    let Vsource1 = V(net1)[i]
    let Vbody1 = V(body1)[i]
    let Id1 = I(Vd)[i]
    let Ig1 = I(Vg1)[i]
    let Is1 = I(Vd2)[i]
    let Ib1 = I(Vb1)[i]
    let Vdrain2 = V(net2)[i]
    let Vgate2 = V(gate2)[i]
    let Vsource2 = V(source2)[i]
    let Vbody2 = V(body2)[i]
    let Id2 = I(Vd2)[i]
    let Ig2 = I(Vg2)[i]
    let Is2 = I(Vs2)[i]
    let Ib2 = I(Vb2)[i]
    echo "$&Vdrain1 $&Vgate1 $&Vsource1 $&Vbody1 $&Id1 $&Ig1 $&Is1 $&Ib1 $&Vdrain2 $&Vgate2 $&Vsource2 $&Vbody2 $&Id2 $&Ig2 $&Is2 $&Ib2" >> NMOS_Stack_00_W1.txt
    let i = i + 1
end

print V(drain1) V(gate1) V(net1) V(body1) I(Vd) I(Vg1) I(Vd2) I(Vb1) V(net2) V(gate2) V(net2) V(body2) I(Vd2) I(Vg2) I(Vs2) I(Vb2)
*end
.ENDC

.END
